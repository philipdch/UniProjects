library verilog;
use verilog.vl_types.all;
entity Exercise_2_vlg_vec_tst is
end Exercise_2_vlg_vec_tst;
