library verilog;
use verilog.vl_types.all;
entity Exercise_2_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exercise_2_vlg_check_tst;
