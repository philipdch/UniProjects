library verilog;
use verilog.vl_types.all;
entity Exercise_1_vlg_sample_tst is
    port(
        X1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic;
        X4              : in     vl_logic;
        X5              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Exercise_1_vlg_sample_tst;
