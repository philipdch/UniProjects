library verilog;
use verilog.vl_types.all;
entity Exercise_3_vlg_vec_tst is
end Exercise_3_vlg_vec_tst;
