library verilog;
use verilog.vl_types.all;
entity Exercise_1_vlg_vec_tst is
end Exercise_1_vlg_vec_tst;
