library verilog;
use verilog.vl_types.all;
entity Exercise_2 is
    port(
        F               : out    vl_logic;
        x2              : in     vl_logic;
        X1              : in     vl_logic;
        x4              : in     vl_logic;
        x3              : in     vl_logic
    );
end Exercise_2;
