library verilog;
use verilog.vl_types.all;
entity ALU_16_Bit_vlg_vec_tst is
end ALU_16_Bit_vlg_vec_tst;
