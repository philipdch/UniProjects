library verilog;
use verilog.vl_types.all;
entity Exercise_3 is
    port(
        X1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic;
        F               : out    vl_logic
    );
end Exercise_3;
